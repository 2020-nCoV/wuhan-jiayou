module main;
  initial
    begin
      $display("💖武汉加油，中国加油🇨🇳!");
      $finish;
    end
endmodule
